module cand
  (
   input       a,b,
   output wire y
   );
   assign y = a & b;
endmodule
